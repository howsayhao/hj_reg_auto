`ifndef __root_map_vh__
`define __root_map_vh__
//**************************************Address Definition Here***************************************//
`define root_map_map_1_TEM21 64'hc//external
`define root_map_map_1_TEM22 64'h10//external
`define root_map_map_1_TEM23 64'h14//external
`define root_map_map_1_TEM21_alias 64'h10c//external
`define root_map_map_1_TEM22_alias 64'h110//external
`define root_map_map_1_TEM23_alias 64'h114//external
`define root_map_shared_map_map_2_shared_2 64'h118//external
`define root_map_shared_map_map_3_shared_3 64'h11c//external
`define root_map_ipxact_map_reg1 64'h200//external
`define root_map_ipxact_map_reg_array0 64'h300//external
`define root_map_ipxact_map_reg_array1 64'h304//external
`define root_map_ipxact_map_reg_array2 64'h308//external
`define root_map_ipxact_map_reg_array3 64'h30c//external
`endif