`ifndef __root_map__root_map__shared_map_vh__
`define __root_map__root_map__shared_map_vh__
//**************************************Address Definition Here***************************************//
`define map_2_shared_2 64'h0//internal
`define map_3_shared_3 64'h4//internal
`endif