`ifndef __test_map_vh__
`define __test_map_vh__
//*************Address Definition Here**************//
`define `test_map_1_inst_test1_TEM21 64'hc//internal
`define `test_map_1_inst_test1_TEM22 64'h10//internal
`define `test_map_1_inst_test1_TEM23 64'h14//internal
`define `test_map_1_inst_test1_TEM21_alias 64'h10c//internal
`define `test_map_1_inst_test1_TEM22_alias 64'h110//internal
`define `test_map_1_inst_test1_TEM23_alias 64'h114//internal
`define `test_map_2_inst_shared_2 64'h118//internal
`define `test_map_3_inst_shared_3 64'h11c//internal
`endif