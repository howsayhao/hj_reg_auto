`ifndef __root_map_vh__
`define __root_map_vh__
//**************************************Address Definition Here***************************************//
`define test_map_2_inst_shared_2 64'h118//internal
`define test_map_3_inst_shared_3 64'h11c//internal
`define reg_t 64'h310//internal
`define test_map_1_inst_TEM21 64'hc//external
`define test_map_1_inst_TEM22 64'h10//external
`define test_map_1_inst_TEM23 64'h14//external
`define test_map_1_inst_TEM21_alias 64'h10c//external
`define test_map_1_inst_TEM22_alias 64'h110//external
`define test_map_1_inst_TEM23_alias 64'h114//external
`define ipxact_block_example_inst_reg1 64'h200//external
`define ipxact_block_example_inst_reg_array0 64'h300//external
`define ipxact_block_example_inst_reg_array1 64'h304//external
`define ipxact_block_example_inst_reg_array2 64'h308//external
`define ipxact_block_example_inst_reg_array3 64'h30c//external
`endif