`ifndef __root_map_vh__
`define __root_map_vh__
//**************************************Address Definition Here***************************************//
`define err_log_0__snap_0 64'h0//internal
`define err_log_0__snap_1 64'h4//internal
`define err_log_1 64'h8//internal
`define root_map_map_1_TEM21 64'h40c//external
`define root_map_map_1_TEM22 64'h410//external
`define root_map_map_1_TEM23 64'h414//external
`define root_map_map_1_TEM21_alias 64'h50c//external
`define root_map_map_1_TEM22_alias 64'h510//external
`define root_map_map_1_TEM23_alias 64'h514//external
`define root_map_shared_map_map_2_shared_2 64'h518//external
`define root_map_shared_map_map_3_shared_3 64'h51c//external
`define root_map_ipxact_map_reg1 64'h600//external
`define root_map_ipxact_map_reg_array0 64'h700//external
`define root_map_ipxact_map_reg_array1 64'h704//external
`define root_map_ipxact_map_reg_array2 64'h708//external
`define root_map_ipxact_map_reg_array3 64'h70c//external
`endif