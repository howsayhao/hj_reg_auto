`ifndef __basic_vh__
`define __basic_vh__
//*************Address Definition Here**************//
`define `foo_r1 64'h0//internal
`define `foo_r2 64'h4//internal
`define `foo_r3 64'h8//internal
`define `bar0_0_r10 64'h1000//internal
`define `bar0_0_r11 64'h1004//internal
`define `bar0_0_r12 64'h1008//internal
`define `bar0_0_r13 64'h100c//internal
`define `bar0_1_r10 64'h1100//internal
`define `bar0_1_r11 64'h1104//internal
`define `bar0_1_r12 64'h1108//internal
`define `bar0_1_r13 64'h110c//internal
`define `bar0_2_r10 64'h1200//internal
`define `bar0_2_r11 64'h1204//internal
`define `bar0_2_r12 64'h1208//internal
`define `bar0_2_r13 64'h120c//internal
`define `bar1_0_r10 64'h1300//internal
`define `bar1_0_r11 64'h1304//internal
`define `bar1_0_r12 64'h1308//internal
`define `bar1_0_r13 64'h130c//internal
`define `bar1_1_r10 64'h1400//internal
`define `bar1_1_r11 64'h1404//internal
`define `bar1_1_r12 64'h1408//internal
`define `bar1_1_r13 64'h140c//internal
`define `bar1_2_r10 64'h1500//internal
`define `bar1_2_r11 64'h1504//internal
`define `bar1_2_r12 64'h1508//internal
`define `bar1_2_r13 64'h150c//internal
`define `bar2_0_r10 64'h1600//internal
`define `bar2_0_r11 64'h1604//internal
`define `bar2_0_r12 64'h1608//internal
`define `bar2_0_r13 64'h160c//internal
`define `bar2_1_r10 64'h1700//internal
`define `bar2_1_r11 64'h1704//internal
`define `bar2_1_r12 64'h1708//internal
`define `bar2_1_r13 64'h170c//internal
`define `bar2_2_r10 64'h1800//internal
`define `bar2_2_r11 64'h1804//internal
`define `bar2_2_r12 64'h1808//internal
`define `bar2_2_r13 64'h180c//internal
`define `bar3_0_r10 64'h1900//internal
`define `bar3_0_r11 64'h1904//internal
`define `bar3_0_r12 64'h1908//internal
`define `bar3_0_r13 64'h190c//internal
`define `bar3_1_r10 64'h1a00//internal
`define `bar3_1_r11 64'h1a04//internal
`define `bar3_1_r12 64'h1a08//internal
`define `bar3_1_r13 64'h1a0c//internal
`define `bar3_2_r10 64'h1b00//internal
`define `bar3_2_r11 64'h1b04//internal
`define `bar3_2_r12 64'h1b08//internal
`define `bar3_2_r13 64'h1b0c//internal
`define `bar2_r10 64'h8000//internal
`define `bar2_r11 64'h8004//internal
`define `bar2_r12 64'h8008//internal
`define `bar2_r13 64'h800c//internal
`define `xxx_r10 64'h10000//external
`define `xxx_r11 64'h10004//external
`define `xxx_r12 64'h10008//external
`define `xxx_r13 64'h1000c//external
`define `xxx_r14 64'h10010//external
`define `xxx_r15 64'h10014//external
`define `xxx_r16 64'h10018//external
`define `xxx_r17 64'h1001c//external
`endif