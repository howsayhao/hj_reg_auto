`ifndef __root_map__root_map__map_1_vh__
`define __root_map__root_map__map_1_vh__
//**************************************Address Definition Here***************************************//
`define TEM21 64'hc//internal
`define TEM22 64'h10//internal
`define TEM23 64'h14//internal
`define TEM21_alias 64'h10c//internal
`define TEM22_alias 64'h110//internal
`define TEM23_alias 64'h114//internal
`endif